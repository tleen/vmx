module vmx

fn init() int {
	println('init called')
	return 1
}

pub fn hello() {
	println('Hello World !')
}
