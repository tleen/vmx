module vmx

fn init() {
	println('init called')
}

pub fn hello() {
	println('Hello World !')
}
