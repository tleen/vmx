module main

import tleen.vmx

fn main() {
	vmx.hello()
}
